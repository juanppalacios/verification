-- log package

-- modeled after Python's logging library: https://docs.python.org/3/library/logging.html

package log_pkg is
    
    type log_level is (none, debug, info, warning, error);
    
    -- log object
    
    
end package;

package body log_pkg is
    
end package body;