-- log package testbench